`timescale 1ns/10ps
module IOTDF( clk, rst, in_en, iot_in, fn_sel, busy, valid, iot_out);
input          clk;
input          rst;
input          in_en;
input  [7:0]   iot_in;
input  [2:0]   fn_sel;
output         busy;
output         valid;
output [127:0] iot_out;

    localparam S_IDLE = 0;
    localparam S_LOAD = 1;
    localparam S_SORT = 2;
    localparam S_DONE = 3;

endmodule
